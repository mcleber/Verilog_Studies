`timescale 1ns / 1ps

module hello_world();

    initial begin
        $display("\n\t Hello World \n");
    end 


endmodule
